//////////////////////////////////////
// ACE GENERATED VERILOG INCLUDE FILE
// Generated on: 2023.06.12 at 14:46:13 PDT
// By: ACE 9.0.1
// From project: vp_project
//////////////////////////////////////
// User Design Port List Include File
//////////////////////////////////////

    // Ports for ethernet_0
    // Clocks and Resets
    input wire        ethernet_0_m0_ff_clk_divby2,
    input wire        ethernet_0_m1_ff_clk_divby2,
    input wire        ethernet_0_ref_clk_divby2,
    // Quad MAC 0 Flow Control
    input wire  [3:0] ethernet_0_quad0_emac_enable,
    input wire  [3:0] ethernet_0_quad0_emac_pause_en,
    input wire  [31:0] ethernet_0_quad0_emac_pause_on,
    output wire [31:0] ethernet_0_quad0_emac_xoff_gen,
    output wire [3:0] ethernet_0_quad0_lpi_txhold,
    output wire [3:0] ethernet_0_quad0_mac_stop_tx,
    output wire [3:0] ethernet_0_quad0_tx_hold_req,
    // Quad MAC 0 Status
    input wire  [3:0] ethernet_0_m0_ffe_tx_ovr,
    input wire  [3:0] ethernet_0_m0_ffp_tx_ovr,
    input wire  [3:0] ethernet_0_m0_mac_tx_underflow,
    // Ports for ethernet_1
    // Clocks and Resets
    input wire        ethernet_1_m0_ff_clk_divby2,
    input wire        ethernet_1_m1_ff_clk_divby2,
    input wire        ethernet_1_ref_clk_divby2,
    // Quad MAC 0 Flow Control
    input wire  [3:0] ethernet_1_quad0_emac_enable,
    input wire  [3:0] ethernet_1_quad0_emac_pause_en,
    input wire  [31:0] ethernet_1_quad0_emac_pause_on,
    output wire [31:0] ethernet_1_quad0_emac_xoff_gen,
    output wire [3:0] ethernet_1_quad0_lpi_txhold,
    output wire [3:0] ethernet_1_quad0_mac_stop_tx,
    output wire [3:0] ethernet_1_quad0_tx_hold_req,
    // Quad MAC 0 Status
    input wire  [3:0] ethernet_1_m0_ffe_tx_ovr,
    input wire  [3:0] ethernet_1_m0_ffp_tx_ovr,
    input wire  [3:0] ethernet_1_m0_mac_tx_underflow 
    // Ports for noc
    // Ports for pll_ddr
    input wire        pll_ddr_lock,
    // Ports for pll_eth_sys_ne_0
    input wire        pll_eth_sys_ne_0_lock,
    // Ports for pll_eth_usr_ne_3
    input wire        i_eth_clk,
    input wire        pll_eth_usr_ne_3_lock,
    // Ports for pll_gddr_SE
    input wire        pll_gddr_SE_lock,
    // Ports for pll_gddr_SW
    input wire        pll_gddr_SW_lock,
    // Ports for pll_noc_ne_1
    input wire        i_clk,
    input wire        i_eth_ts_clk,
    input wire        i_reg_clk,
    input wire        pll_noc_ne_1_lock,
    // Ports for pll_pcie
    input wire        pll_pcie_lock,
    // Ports for vp_clkio_ne
    input wire        fpga_rst_l,
    // Ports for vp_clkio_nw
    // Ports for vp_clkio_se
    // Ports for vp_clkio_sw
    // Ports for vp_gpio_n_b0
    // Core Data
    // Port name: ext_gpio_fpga_in[0] has been automatically combined into a the bussed signal below.
    input wire        ext_gpio_fpga_in[7:0],
    // Port name: ext_gpio_fpga_in[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[7] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[0] has been automatically combined into a the bussed signal below.
    output wire       ext_gpio_fpga_oe[7:0],
    // Port name: ext_gpio_fpga_oe[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[7] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[0] has been automatically combined into a the bussed signal below.
    output wire       ext_gpio_fpga_out[7:0],
    // Port name: ext_gpio_fpga_out[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[7] has been automatically combined into a bussed signal.
    output wire       ext_gpio_oe_l,
    output wire       ext_gpio_oe_l_oe,
    output wire       led_oe_l,
    output wire       led_oe_l_oe,
    // Ports for vp_gpio_n_b1
    // Core Data
    // Port name: ext_gpio_dir[0] has been automatically combined into a the bussed signal below.
    output wire       ext_gpio_dir[7:0],
    // Port name: ext_gpio_dir[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[7] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[0] has been automatically combined into a the bussed signal below.
    output wire       ext_gpio_dir_oe[7:0],
    // Port name: ext_gpio_dir_oe[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[7] has been automatically combined into a bussed signal.
    // Port name: led_l[4] has been automatically combined into a the bussed signal below.
    output wire       led_l[7:0],
    // Port name: led_l[5] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[4] has been automatically combined into a the bussed signal below.
    output wire       led_l_oe[7:0],
    // Port name: led_l_oe[5] has been automatically combined into a bussed signal.
    // Ports for vp_gpio_n_b2
    // Core Data
    // Port name: led_l[0] has been automatically combined into a bussed signal.
    // Port name: led_l[1] has been automatically combined into a bussed signal.
    // Port name: led_l[2] has been automatically combined into a bussed signal.
    // Port name: led_l[3] has been automatically combined into a bussed signal.
    // Port name: led_l[6] has been automatically combined into a bussed signal.
    // Port name: led_l[7] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[0] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[1] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[2] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[3] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[6] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[7] has been automatically combined into a bussed signal.
    // Ports for vp_gpio_s_b0
    // Core Data
    input wire        fpga_avr_rxd,
    input wire        fpga_ftdi_rxd,
    input wire        fpga_i2c_mux_gnt,
    input wire        irq_to_fpga,
    input wire        qsfp_int_fpga_l,
    output wire       fpga_avr_txd,
    output wire       fpga_avr_txd_oe,
    output wire       fpga_ftdi_txd,
    output wire       fpga_ftdi_txd_oe,
    output wire       fpga_i2c_req_l,
    output wire       fpga_i2c_req_l_oe,
    output wire       irq_to_avr,
    output wire       irq_to_avr_oe,
    // Port name: test[1] has been automatically combined into a the bussed signal below.
    output wire       test[2:1],
    // Port name: test_oe[1] has been automatically combined into a the bussed signal below.
    output wire       test_oe[2:1],
    // Ports for vp_gpio_s_b1
    // Core Clock
    input wire        mcio_vio_45_10_clk,
    // Core Data
    // Port name: mcio_vio_in[0] has been automatically combined into a the bussed signal below.
    input wire        mcio_vio_in[3:0],
    // Port name: mcio_vio_in[1] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_in[2] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_in[3] has been automatically combined into a bussed signal.
    // Port name: mcio_dir[0] has been automatically combined into a the bussed signal below.
    output wire       mcio_dir[3:0],
    // Port name: mcio_dir[1] has been automatically combined into a bussed signal.
    // Port name: mcio_dir[2] has been automatically combined into a bussed signal.
    // Port name: mcio_dir[3] has been automatically combined into a bussed signal.
    output wire       mcio_dir_45,
    output wire       mcio_dir_45_oe,
    // Port name: mcio_dir_oe[0] has been automatically combined into a the bussed signal below.
    output wire       mcio_dir_oe[3:0],
    // Port name: mcio_dir_oe[1] has been automatically combined into a bussed signal.
    // Port name: mcio_dir_oe[2] has been automatically combined into a bussed signal.
    // Port name: mcio_dir_oe[3] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_oe[0] has been automatically combined into a the bussed signal below.
    output wire       mcio_vio_oe[3:0],
    // Port name: mcio_vio_oe[1] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_oe[2] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_oe[3] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_out[0] has been automatically combined into a the bussed signal below.
    output wire       mcio_vio_out[3:0],
    // Port name: mcio_vio_out[1] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_out[2] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_out[3] has been automatically combined into a bussed signal.
    // Port name: test[2] has been automatically combined into a bussed signal.
    // Port name: test_oe[2] has been automatically combined into a bussed signal.
    // Ports for vp_gpio_s_b2
    // Core Data
    input wire        fpga_sys_scl_in,
    input wire        fpga_sys_sda_in,
    input wire        mcio_scl_in,
    input wire        mcio_sda_in,
    output wire       fpga_sys_scl_oe,
    output wire       fpga_sys_scl_out,
    output wire       fpga_sys_sda_oe,
    output wire       fpga_sys_sda_out,
    output wire       mcio_oe1_l,
    output wire       mcio_oe1_l_oe,
    output wire       mcio_oe_45_l,
    output wire       mcio_oe_45_l_oe,
    output wire       mcio_scl_oe,
    output wire       mcio_scl_out,
    output wire       mcio_sda_oe,
    output wire       mcio_sda_out,
    // Ports for vp_pll_nw_2
    input wire        pll_nw_2_ref0_312p5_clk,
    input wire        vp_pll_nw_2_lock,
    // Ports for vp_pll_sw_2
    input wire        pll_sw_2_ref1_312p5_clk,
    input wire        vp_pll_sw_2_lock,

//////////////////////////////////////
// End User Design Port List Include File
//////////////////////////////////////
